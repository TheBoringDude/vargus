module vargus

