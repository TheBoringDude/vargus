module vargus

fn (v &Vargus) help() {
	
}