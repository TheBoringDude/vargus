module vargus

pub fn (c &Commander) help() {
	println(c)
}